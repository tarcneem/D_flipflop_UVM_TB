
`ifndef DFF_INTF_SV
`define DFF_INTF_SV
interface dff_intf;
    logic clk;
    logic rst;
    logic din;
    logic dout;
  endinterface
`endif