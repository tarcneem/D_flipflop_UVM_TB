`include "dff_intf.sv"
`include "sequence_item.sv"
`include "sequence_dff.sv"
`include "sequencer.sv"
`include "driver_dff.sv"
`include "monitor_dff.sv"
`include "agent_dff.sv"
`include "scoreboard_dff.sv"
`include "Env.sv"
`include "test_dff.sv"
