import uvm_pkg::*;
`include "uvm_macros.svh"
`include "sequence_item.sv" 
`ifndef SEQUENCER_SV
`define SEQUENCER_SV
class sequencer extends uvm_sequencer#(sequence_item);
`uvm_component_utils(sequencer)

    function new(string name="sequencer",uvm_component parent);
        super.new(name,parent);
    endfunction
endclass
`endif